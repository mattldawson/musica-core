netcdf chebev_coeffs {
dimensions:
	nchebev_wave = 17 ;
  nchebev_wave_edge = 18 ;
	nchebev_term = 20 ;
variables:
  double wl_edge(nchebev_wave_edge) ;
    wl_edge:description = "wavelength edge" ;
    wl_edge:units = "nm" ;
    wl_edge:long_name = "wavelength edge" ;
	double chebev_ac(nchebev_wave, nchebev_term) ;
		chebev_ac:description = "chebev a coefficient" ;
		chebev_ac:units = "none" ;
		chebev_ac:longname = "chebev a coefficient" ;
	double chebev_bc(nchebev_wave, nchebev_term) ;
		chebev_bc:description = "chebev b coefficient" ;
		chebev_bc:units = "none" ;
		chebev_bc:longname = "chebev b coefficient" ;

// global attributes:
		:history = "Wed Jul 10 13:30:26 2019: ncks -v chebev_ac,chebev_bc wrf_tuv_xsqy.nc chebev_coeffs.nc" ;
		:NCO = "netCDF Operators version 4.7.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 wl_edge =
   174.4, 177.0, 178.6, 180.2, 181.8, 183.5, 185.2, 186.9, 188.7,
   190.5, 192.3, 194.2, 196.1, 198.0, 200.0, 202.0, 204.1, 205.8 ;

 chebev_ac =
  0.0101299248635769, 0.00492775812745094, -0.00321849016472697, 
    -0.00222120410762727, -0.0011063467245549, -0.000602349755354226, 
    -0.00053768081124872, -0.000352014612872154, -9.80006880126894e-05, 
    0.000391476933145896, 0.000375378964236006, -4.47879792773165e-05, 
    -8.38850537547842e-05, 7.58726091589779e-05, 5.0431837735232e-05, 
    -0.000130119049572386, -0.000133143141283654, 8.9079316239804e-05, 
    6.90536253387108e-05, -0.000112801055365708,
  0.0124629074707627, 0.00669141532853246, -0.00361971813254058, 
    -0.00454070419073105, -0.00308012403547764, -0.000475269422167912, 
    -0.000122243043733761, -0.000409653090173379, -0.000166980593348853, 
    0.0001743208267726, 0.000428983476012945, 0.000358218618202955, 
    -0.000190981372725219, -0.000211607097298838, 0.000290705938823521, 
    2.1953013856546e-05, -0.000401182536734268, -3.48842986568343e-05, 
    0.000211630875128321, 5.28662712895311e-06,
  0.0117507819086313, 0.00674931425601244, -0.00171727291308343, 
    -0.00243034074082971, -0.00169446307700127, 0.000154578810906969, 
    0.000568136456422508, 0.000364597071893513, -0.000206275508389808, 
    -0.000553898862563074, 4.62679454358295e-05, 0.00048778869677335, 
    -2.66857368842466e-05, -0.000299255974823609, 0.000142124335980043, 
    0.000101043260656297, -0.000206791257369332, 7.05252678017132e-05, 
    0.000131553868413903, -0.00018564480706118,
  0.00600254954770207, 0.00304163340479136, -0.00134564808104187, 
    -3.05988360196352e-05, 0.000544505892321467, 2.08055030270771e-06, 
    -7.8972960182e-05, 0.000369826360838488, 7.07908038748428e-05, 
    -0.000194968146388419, -0.000145655474625528, -9.36690485104918e-05, 
    8.34015081636608e-05, 0.000131876877276227, 2.86733734355948e-06, 
    -5.55848673684523e-05, -6.40066064079292e-05, -1.81727118615527e-05, 
    7.14663256076165e-05, 7.83157447585836e-05,
  0.00383285153657198, 0.00092475104611367, -0.00241587474010885, 
    -0.000750405946746469, 0.000121707023936324, -4.61681847809814e-05, 
    -0.000261324108578265, 1.65143301273929e-05, -4.79382542835083e-05, 
    -0.000120529599371366, -1.09635375338257e-05, 2.28264107136056e-05, 
    5.02281145600136e-05, 8.85566769284196e-05, 5.17402586410753e-05, 
    -0.000105991442978848, -0.000150590596604161, 6.29041242063977e-05, 
    0.000126962651847862, -2.21114532905631e-05,
  0.00419552065432072, -6.93289621267468e-05, -0.00142452772706747, 
    -0.000860366330016404, 0.000208176628802903, -0.000203694653464481, 
    -0.000458434136817232, 9.22639737837017e-05, 0.000148562714457512, 
    -9.61433397606015e-05, -0.000165128527441993, -5.45398215763271e-05, 
    0.000123535690363497, 0.000169545091921464, 4.28201747126877e-05, 
    -0.000132499873870984, -0.000165795601787977, 1.55489578901324e-05, 
    0.000140164876938798, 6.84259503032081e-05,
  0.0086836451664567, 0.00365910609252751, 0.000817305641248822, 
    0.000605895183980465, 0.00135609519202262, 0.000594568497035652, 
    -0.000300284940749407, -0.000462242780486122, -0.000473478634376079, 
    -0.000247934163780883, -8.93372707650997e-05, -0.000107828869658988, 
    0.000123617821373045, 0.000366481574019417, 0.000207662509637885, 
    -0.000137203343911096, -0.000318799575325102, -0.000172551663126796, 
    0.000198595487745479, 0.000331698509398848,
  0.00661816960200667, -0.000216037646168843, 0.000140400865348056, 
    -0.00117858254816383, 0.000611105002462864, -5.91504394833464e-05, 
    -0.000630654161795974, -6.64311737637036e-05, -5.13576233061031e-05, 
    -0.000101171179267112, -0.000179289738298394, -0.000205253978492692, 
    0.000120076554594561, 0.000339650665409863, 0.000141964104841463, 
    -9.84250364126638e-05, -0.000210368321859278, -0.000165707358974032, 
    0.000117976356705185, 0.000260581320617348,
  0.00545611511915922, -0.00362338265404105, -0.00136525114066899, 
    -0.00360865192487836, -0.000619182654190809, -0.000434186658822, 
    -0.000804820447228849, -0.00027433640207164, -0.000156403053551912, 
    6.0632035456365e-05, 2.66725837718695e-05, -6.46504267933778e-05, 
    0.000136898175696842, 0.000258964777458459, 8.20863861008547e-05, 
    -0.000166028941748664, -0.000286052090814337, -0.000116959294246044, 
    0.000226951873628423, 0.00027232023421675,
  0.00937877129763365, -0.00100316479802132, -0.00031705157016404, 
    -0.000608240137808025, 0.000772952742408961, 0.000381475576432422, 
    0.000525643583387136, 0.000368972570868209, -0.000559872714802623, 
    -0.000548409123439342, -0.000169998835190199, -1.51356452988693e-05, 
    0.0001343603071291, 0.000216271728277206, 0.000160308176418766, 
    -4.6649387513753e-05, -0.000266584218479693, -0.000129552005091682, 
    0.000200681111891754, 0.000218566958210431,
  0.003731933189556, -0.00214893510565162, -0.00124988087918609, 
    -0.00427354173734784, -0.00169471651315689, -0.00078980007674545, 
    -0.00056980864610523, -0.000137156908749603, -0.000171511404914781, 
    2.2579441065318e-05, -3.77506330551114e-05, -0.000183850948815234, 
    4.12766639783513e-05, 0.000240967245190404, 0.000104495644336566, 
    -0.000112460977106821, -0.000205384247237816, -8.39542481116951e-05, 
    0.000187522658961825, 0.000233914193813689,
  0.00425203470513225, -0.00402387976646423, 0.000252219004323706, 
    -0.00403935508802533, -0.000614812306594104, -5.09671117470134e-05, 
    -0.000203741161385551, 1.97204317373689e-05, -0.000450919003924355, 
    -0.000126005616039038, 8.93721517059021e-05, -2.71678818535293e-05, 
    5.80054256715812e-05, 0.000130286993226036, 3.37692035827786e-05, 
    -3.93697191611864e-05, -0.000101442463346757, -8.10016208561137e-05, 
    9.08265137695707e-05, 0.000107638246845454,
  0.0111884698271751, -0.00815672241151333, 0.00505659403279424, 
    -0.00570040382444859, 0.00100072589702904, 0.000859443447552621, 
    -9.43752093007788e-06, 0.000551758916117251, -0.000782699382398278, 
    -0.00028945694793947, 0.000196798151591793, -1.76409503183095e-05, 
    2.83752870018361e-05, 5.05548741784878e-05, -5.16218606207985e-05, 
    2.88155551970704e-05, -3.08373643065352e-07, -6.93029578542337e-05, 
    8.83697211975232e-05, 2.91644864773843e-05,
  0.0122261606156826, -0.00848923996090889, 0.00496717588976026, 
    -0.00458617974072695, 0.000975968316197395, 0.000716903537977487, 
    -0.000238989494391717, 0.000550234690308571, -0.000412657798733562, 
    -0.000235748302657157, 4.87558972963598e-05, -8.5518098785542e-05, 
    1.29317804749007e-05, 8.10621932032518e-05, -1.54078370542265e-05, 
    2.44258608290693e-05, 1.30732860270655e-05, -6.1198414186947e-05, 
    4.75925880891737e-05, 1.97788322111592e-05,
  0.00658877100795507, -0.00433475291356444, 0.00263612275011837, 
    -0.00221549510024488, 0.00068632181501016, 0.000227582058869302, 
    -0.00012734139454551, 0.000365001847967505, -0.000265894341282547, 
    -0.000130875501781702, 4.99247180414386e-05, -3.80796154786367e-05, 
    1.90326791198459e-05, 2.66042261500843e-05, -2.8188720534672e-05, 
    3.08026319544297e-05, 1.63951899594394e-05, -4.17931187257636e-05, 
    2.42550577240763e-05, 5.66097878618166e-06,
  0.0021509004291147, -0.00166029925458133, 0.00118536711670458, 
    -0.000912618008442223, 0.000250681827310473, 8.15023668110371e-05, 
    -7.89691766840406e-05, 0.000130603119032457, -0.000102240068372339, 
    -4.33807872468606e-05, 2.61714540101821e-05, -1.57990307343425e-05, 
    2.62594153355167e-06, 9.48948127188487e-06, -1.00102888609399e-05, 
    1.39703633976751e-05, 9.96544440567959e-06, -1.6860552932485e-05, 
    5.0446665227355e-06, -1.07585015030054e-06,
  0.000719559495337307, -0.000414013979025185, 0.000426325888838619, 
    -0.000208456083782949, 0.00011891005851794, 6.36485347058624e-05, 
    -1.1551941270227e-06, 4.96710745210294e-05, -2.94810397463152e-05, 
    -2.04631523956778e-05, 4.90748880110914e-06, -5.67996175959706e-06, 
    -2.67588825408893e-06, 1.94920335161441e-06, -1.04792957245081e-06, 
    5.66770722798537e-06, 4.32715751230717e-06, -4.63129254058003e-06, 
    4.18031902427174e-07, -4.08798939588451e-07 ;

 chebev_bc =
  -90.3405380249023, -2.04607248306274, 0.551205933094025, 0.260696977376938, 
    -0.193879470229149, -0.0922096222639084, 0.100352182984352, 
    0.00635678973048925, -0.021759707480669, -0.0289956964552402, 
    0.0162216145545244, 0.0204767286777496, -0.0173658542335033, 
    -0.00330401235260069, 0.0115237347781658, -0.00141748634632677, 
    -0.00472612958401442, 0.00052261893870309, 0.00113617908209562, 
    -0.0010145918931812,
  -93.2331466674805, -3.16542029380798, 0.6362424492836, 0.39213439822197, 
    -0.144075363874435, -0.0932125896215439, 0.0178563371300697, 
    -0.0104700718075037, 0.029554920271039, -0.0189487375319004, 
    -0.00735823297873139, 0.0138181876391172, -0.00441416772082448, 
    0.000395223614759743, 0.00129860453307629, -0.00456838915124536, 
    0.00284727034159005, 0.00898296944797039, -0.00268963188864291, 
    -0.015950683504343,
  -93.8624114990234, -2.94678354263306, 0.578123450279236, 0.388009339570999, 
    -0.146021634340286, -0.070644348859787, 0.0450663156807423, 
    -0.0511583872139454, 0.0261675920337439, 0.0182473622262478, 
    -0.0120020741596818, 0.00589253241196275, -0.0109326224774122, 
    -0.00778053374961019, 0.0153118809685111, 0.00407321099191904, 
    -0.0105885416269302, 0.000580691616050899, 0.00559028051793575, 
    -0.00530823273584247,
  -94.0979385375977, -2.90637922286987, 0.353586196899414, 0.55381977558136, 
    -0.117143325507641, -0.141220405697823, 0.0482261255383492, 
    -0.0235740207135677, 0.0202542319893837, 0.028289046138525, 
    -0.017188360914588, -0.0134796556085348, 0.00362913589924574, 
    0.00382174691185355, 0.000842229928821325, 2.48882333835354e-05, 
    -0.000953577051404864, 0.000493692758027464, 0.000750306702684611, 
    -0.00248248502612114,
  -95.3380661010742, -3.08791637420654, 0.275621891021729, 0.57646244764328, 
    -0.0762977302074432, -0.142043337225914, 0.0323133505880833, 
    -0.0209645349532366, 0.0173386912792921, 0.0159379933029413, 
    -0.0151440035551786, 0.00195670663379133, 0.00524273794144392, 
    -0.00828419532626867, -0.00236440217122436, 0.00531308772042394, 
    0.00231126416474581, 0.0023872833698988, -0.00132964784279466, 
    -0.00878510251641273,
  -96.4176712036133, -2.85797882080078, 0.0582633949816227, 
    0.637516021728516, -0.05312330275774, -0.148185417056084, 
    0.0288811642676592, -0.0107717551290989, -0.0111621981486678, 
    0.0298001021146774, 0.00823272950947285, -0.0183217860758305, 
    -0.00245161238126457, 0.00180326553527266, -0.00395141821354628, 
    0.00607215240597725, 0.00678080320358276, -0.00374749070033431, 
    -0.00499235698953271, -0.000664978986606002,
  -97.0311737060547, -2.59352040290833, -0.0702516734600067, 
    0.600104868412018, 0.015121947042644, -0.163790091872215, 
    0.00744506483897567, 0.0109807569533587, -0.0219006221741438, 
    0.0175820365548134, 0.0266449004411697, -0.012944795191288, 
    -0.0187923610210419, -0.0018237226177007, 0.00182844023220241, 
    0.0072054285556078, 0.0103801088407636, -0.000637304387055337, 
    -0.00960146356374025, -0.00667825061827898,
  -98.6436004638672, -2.53565645217896, -0.329384177923203, 
    0.650445640087128, 0.0522664524614811, -0.105886295437813, 
    -0.0272549111396074, 0.014848162420094, -0.0013233054196462, 
    0.000113022615551017, 0.0175962075591087, -0.0101386746391654, 
    -0.00908265728503466, 0.001663449103944, -0.00244091334752738, 
    0.00407648412510753, 0.0088880667462945, 0.000557112856768072, 
    -0.00829594302922487, -0.00501646054908633,
  -100.008163452148, -2.25186800956726, -0.515524744987488, 
    0.624725878238678, 0.0604026541113853, -0.0832023620605469, 
    -0.0638432949781418, 0.0168268624693155, -0.0072116032242775, 
    -0.0222005303949118, 0.0361178927123547, 0.0107328006997705, 
    -0.0176986623555422, -0.0130304899066687, -0.000123355697724037, 
    0.00989387370646, 0.00833328813314438, 0.00349754258058965, 
    -0.00898257363587618, -0.0119734387844801,
  -101.109031677246, -2.08251047134399, -0.485277205705643, 
    0.480242609977722, 0.135131850838661, -0.0687109902501106, 
    -0.0555102564394474, 0.0311791598796844, 0.00463733728975058, 
    -0.017877385020256, 0.0227369107306004, 0.00596637604758143, 
    -0.0176265612244606, -0.0113650029525161, 0.00496777752414346, 
    0.011115426197648, 0.00327587174251676, -0.000773543084505945, 
    -0.00497137242928147, -0.00657283561304212,
  -101.378021240234, -2.06618666648865, -0.750329852104187, 
    0.474477708339691, 0.216930583119392, -0.00205568270757794, 
    -0.136293798685074, -0.0208189357072115, 0.0336209423840046, 
    -0.0095396526157856, 0.00507326703518629, 0.00816291105002165, 
    0.00254143308848143, -0.0126592088490725, -0.0124136367812753, 
    0.00966589339077473, 0.0146281374618411, 0.00240311096422374, 
    -0.0106695694848895, -0.00910557806491852,
  -102.960906982422, -1.33756220340729, -0.749491631984711, 
    0.420921385288239, 0.0905516892671585, 0.0524549372494221, 
    -0.128325313329697, -0.0217408537864685, 0.0523338168859482, 
    -0.00580802280455828, -0.00191919889766723, -0.0115864919498563, 
    0.00611819559708238, 0.00531047722324729, -0.00836107321083546, 
    0.000184082484338433, 0.00508535699918866, 0.00462298654019833, 
    -0.00460129836574197, -0.00562931969761848,
  -105.169540405273, -0.205385372042656, -0.918219983577728, 
    0.64212566614151, -0.200856730341911, 0.173608526587486, 
    -0.139732763171196, -0.0203941967338324, 0.0747282952070236, 
    -0.0288790408521891, 0.0184939019382, -0.0248577445745468, 
    0.00110148615203798, 0.0127701479941607, -0.00647783745080233, 
    0.00191333214752376, -0.00258093187585473, 0.00393378455191851, 
    -0.00175894307903945, -0.000816778454463929,
  -106.506790161133, 0.391759157180786, -0.67700332403183, 0.452103555202484, 
    -0.257609605789185, 0.186408057808876, -0.0743092522025108, 
    -0.0268692187964916, 0.0396465323865414, -0.0295525956898928, 
    0.0294464193284512, -0.0123819792643189, -0.00574772898107767, 
    0.00414400268346071, -0.00401446921750903, 0.00559650314971805, 
    -0.00148067332338542, 0.000972851878032088, -0.00207512849010527, 
    0.000830528151709586,
  -106.438453674316, 0.196900457143784, -0.380969196557999, 0.24158650636673, 
    -0.13838629424572, 0.103819482028484, -0.0392660833895206, 
    -0.0125685445964336, 0.0188454631716013, -0.0177583992481232, 
    0.0179644040763378, -0.00642563076689839, -0.00294574745930731, 
    0.00203659082762897, -0.00275633274577558, 0.00334151485003531, 
    -0.000784205738455057, 0.00038380260230042, -0.00103575247339904, 
    0.000640276586636901,
  -106.576293945313, 0.114275127649307, -0.142852753400803, 
    0.0971360057592392, -0.0631433874368668, 0.04073765873909, 
    -0.013855554163456, -0.00303270015865564, 0.00803583581000566, 
    -0.0086203096434474, 0.0060861399397254, -0.00250944681465626, 
    -0.000381184683647007, 0.00142290280200541, -0.00120228028390557, 
    0.000858944142237306, -0.000630583963356912, 0.000224662348045968, 
    -0.00014879037917126, 0.000516644853632897,
  -106.590606689453, 0.0423569343984127, -0.0367124788463116, 
    0.0293931346386671, -0.0193247962743044, 0.0106352576985955, 
    -0.00423215143382549, -0.000530433084350079, 0.00294468132779002, 
    -0.00227004685439169, 0.0016710382187739, -0.000828482676297426, 
    -0.00030543448519893, 0.000429603038355708, -0.000243537855567411, 
    0.000240759894950315, -0.000196340362890624, 4.22856719524134e-05, 
    -2.52488480327884e-05, 0.000172790678334422 ;
}
